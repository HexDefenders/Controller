`timescale 1ns / 1ps

module glyphs #(parameter WIDTH = 64, ADR_BITS = 8) 
				   (clk, en, value, glyph);
	input clk, en;
	input [ADR_BITS-1:0] value;
	output reg [WIDTH-1:0] glyph;
	
	reg [WIDTH-1:0] glyphs [(2*ADR_BITS)-1:0];
	
	initial begin
	
		// To generate other glyphs: http://robojax.com/learn/arduino/8x8LED/
		// NOTE: reverse the order of each row (column: right to left, row: top to bottom)
		glyphs[8'h0] = 64'b0000000000011100001000100010001000100010001000100010001000011100;
		glyphs[8'h1] = 64'b0000000000000100000001000000011000000110000001100000011000000110;
		glyphs[8'h2] = 64'b0000000000001100000100100001000000001000000001000000001000011110;
		glyphs[8'h3] = 64'b0000000000011100001000100010000000011000001000000010001000011100;
		glyphs[8'h4] = 64'b0000000000100010001000100010001000111110001000000010000000100000;
		glyphs[8'h5] = 64'b0000000000111110000000100000001000011110001000000010000000011110;
		glyphs[8'h6] = 64'b0000000000011100000000100000001000011010001001100010001000011100;
		glyphs[8'h7] = 64'b0000000000011110000100000001000000111100000010000000010000000010;
		glyphs[8'h8] = 64'b0000000000011100001000100010001000011100001000100010001000011100;
		glyphs[8'h9] = 64'b0000000000011100001000100010001000111100001000000010001000011100;
		glyphs[8'ha] = 64'b0000000000011000001001000100001001000010011111100100001001000010;
		glyphs[8'hb] = 64'b0000000000011110001000100010001000011110001000100010001000011110;
		glyphs[8'hc] = 64'b0000000000011000001001000000001000000010000000100010010000011000;
		glyphs[8'hd] = 64'b0000000000001110000100100010001000100010001000100001001000001110;
		glyphs[8'he] = 64'b0000000000111110000000100000001000011110000000100000001000111110;
		glyphs[8'hf] = 64'b0000000000111110000000100000001000011110000000100000001000000010;
//		glyphs[5'h10] = 64'b0000000000000000000000000100010000101000000100000010100001000100; // x
	
	end
	
	always @(posedge clk)
		if (en)
			glyph <= glyphs[value]; 
	
endmodule
